module CRUDE_AWAKENING(
     input wire       in0,
     output wire       out
);
    assign out = in0;
endmodule
