module test_module (
    input    i_data1, // 入力信号線の定義
    input    i_data2,
    output   o_data1  // 出力信号線の定義
);
 // 回路
endmodule