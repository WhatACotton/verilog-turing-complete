module BYTE_NOT(
     input wire [7:0] in0,
     output wire [7:0] out
);

endmodule